//CLASS
`timescale 1n/100ps

//INTERFAZ
        //CLOCKINGBLOCKS Y MODPORTS ESTAN DENTRO DE LA INTERFAZ?
    //CLOCKINGBLOCKS

    //MODPORTS
//ENDINTERFACE

//CLASS SCOREBOARD

//TASK MONITOR INPUT
//TASK MONITOR OUTPUT

//PROGRAM

    //COVERGROUPS
    //DECLARACION OBJETOS Y COVERGROUPS
    //INITIAL
        //CREAMOS LOS OBJETOS
        //LANZAMOS PROCEDIMIENTO

        //WHILES ACTIVACIONES CONSTRAINTS

//ENDPROGAM
module tb_top_aleatorizado (
);
//DECLARACIONES SEÑALES

//INSTANCIACION INTERFAZ

//INSTANCIACION DUV

//LLAMADA A PROGAM

//GENERACIOND EL RELOJ

//INITIAL

endmodule